// `timescale 1ns / 1ps

`include "top.sv"
`include "single_port_ram.sv"